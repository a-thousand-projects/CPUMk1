library verilog;
use verilog.vl_types.all;
entity tb_Mux4x16 is
end tb_Mux4x16;

library verilog;
use verilog.vl_types.all;
entity mux_test is
end mux_test;
